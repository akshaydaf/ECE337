/home/ecegrid/a/mg27/ece337/Lab2/source/tb_adder_1bit.sv