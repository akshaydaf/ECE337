/home/ecegrid/a/mg27/ece337/Lab2/source/adder_8bit.sv